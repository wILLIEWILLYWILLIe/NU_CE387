
`ifndef CORDIC_GLOBAL_SV
`define CORDIC_GLOBAL_SV

parameter string RAD_FILE_NAME = "../source/rad.txt";
parameter string SIN_FILE_NAME = "../source/sin.txt";
parameter string COS_FILE_NAME = "../source/cos.txt";

`endif
