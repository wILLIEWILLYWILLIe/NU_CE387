`ifndef __GLOBALS__
`define __GLOBALS__

// UVM Globals
localparam string PCAP_INPUT_NAME = "../ref/test.pcap";
localparam string REF_OUTPUT_NAME = "../ref/test_output.txt";

`endif
