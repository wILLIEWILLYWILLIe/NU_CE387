
`ifndef CORDIC_SEQUENCE_SV
`define CORDIC_SEQUENCE_SV

class cordic_sequence extends uvm_sequence#(cordic_transaction);
    `uvm_object_utils(cordic_sequence)

    function new(string name = "cordic_sequence");
        super.new(name);
    endfunction

    virtual task body();
        int fd;
        int code;
        logic signed [31:0] rad_val;
        
        // Open the stimulus file (generated by C++ model)
        fd = $fopen(RAD_FILE_NAME, "r");
        if (fd == 0) begin
            `uvm_fatal("SEQ", $sformatf("Could not open %s", RAD_FILE_NAME))
        end

        while (!$feof(fd)) begin
            code = $fscanf(fd, "%h\n", rad_val);
            if (code != 1) break;

            req = cordic_transaction::type_id::create("req");
            start_item(req);
            req.rad_in = rad_val;
            finish_item(req);
        end
        
        $fclose(fd);
    endtask

endclass

`endif
