
module grayscale (
    input  logic        clock,
    input  logic        reset,
    output logic        in_rd_en,
    input  logic        in_empty,
    input  logic [23:0] in_dout,
    output logic        out_wr_en,
    input  logic        out_full,
    output logic [7:0]  out_din
);

    typedef enum logic [0:0] {s0, s1} state_types;
    state_types state, state_c;

    logic [7:0] gs, gs_c;

    always_ff @(posedge clock or posedge reset) begin
        if (reset == 1'b1) begin
            state <= s0;
            gs <= 8'h0;
        end else begin
            state <= state_c;
            gs <= gs_c;
        end
    end

    always_comb begin
        in_rd_en  = 1'b0;
        out_wr_en = 1'b0;
        out_din   = 8'b0;
        state_c   = state;
        gs_c = gs;

        case (state)
            s0: begin
                if (in_empty == 1'b0) begin
                    // Standard division to ensure bit-true accuracy
                    gs_c = 8'(($unsigned({2'b0, in_dout[23:16]}) + $unsigned({2'b0, in_dout[15:8]}) + $unsigned({2'b0, in_dout[7:0]})) / $unsigned(10'd3));
                    in_rd_en = 1'b1;
                    state_c = s1;
                end
            end

            s1: begin
                if (out_full == 1'b0) begin
                    out_din = gs;
                    out_wr_en = 1'b1;
                    state_c = s0;
                end
            end

            default: begin
                in_rd_en  = 1'b0;
                out_wr_en = 1'b0;
                out_din = 8'b0;
                state_c = s0;
                gs_c = 8'hX;
            end

        endcase
    end

endmodule
