
module cordic_tb;

    logic        clock;
    logic        reset;
    logic        valid_in;
    logic signed [31:0] rad_in;
    logic        valid_out;
    logic signed [15:0] sin_out;
    logic signed [15:0] cos_out;

    // File handles and data
    integer rad_file, sin_file, cos_file;
    integer r_scan;
    logic signed [31:0] rad_ref;
    logic signed [15:0] sin_ref;
    logic signed [15:0] cos_ref;
    
    integer errors = 0;
    integer tests = 0;

    // DUT Instance
    logic fifo_full;

    cordic_top dut (
        .clock(clock),
        .reset(reset),
        .valid_in(valid_in),
        .rad_in(rad_in),
        .full_out(fifo_full), // Connect Full
        .valid_out(valid_out),
        .sin_out(sin_out),
        .cos_out(cos_out)
    );

    // Clock Generation
    initial begin
        clock = 0;
        forever #5 clock = ~clock;
    end

    // Cycle Counting
    integer cycle_count = 0;
    integer start_cycle = 0;
    integer latency = 0;
    integer total_latency = 0;
    
    always @(posedge clock) begin
        if (reset) cycle_count <= 0;
        else cycle_count <= cycle_count + 1;
    end

    // Test Procedure
    initial begin
        // Open files (locally generated by C++ model)
        rad_file = $fopen("../source/rad.txt", "r");
        sin_file = $fopen("../source/sin.txt", "r");
        cos_file = $fopen("../source/cos.txt", "r");

        if (rad_file == 0 || sin_file == 0 || cos_file == 0) begin
            $display("Error: Could not open reference files. Run C++ model first.");
            $finish;
        end

        // Reset
        reset = 1;
        valid_in = 0;
        rad_in = 0;
        repeat (5) @(posedge clock);
        reset = 0;
        repeat (5) @(posedge clock);

        // Drive Inputs
        while (!$feof(rad_file) && !$feof(sin_file) && !$feof(cos_file)) begin
            r_scan = $fscanf(rad_file, "%h\n", rad_ref);
            if (r_scan != 1) break; 
            
            // Read expected outputs
            r_scan = $fscanf(sin_file, "%h\n", sin_ref);
            r_scan = $fscanf(cos_file, "%h\n", cos_ref);

            @(posedge clock);
            while (fifo_full) @(posedge clock); // Wait if FIFO is full
            valid_in = 1;
            rad_in = rad_ref;
            start_cycle = cycle_count; // Capture start cycle
            
            @(posedge clock);
            valid_in = 0;

            wait(valid_out);
            latency = cycle_count - start_cycle;
            total_latency = total_latency + latency;
            
            // Check results
            if (sin_out !== sin_ref || cos_out !== cos_ref) begin
                $display("Error at test %0d: rad=%h | exp sin=%h cos=%h | got sin=%h cos=%h", 
                         tests, rad_ref, sin_ref, cos_ref, sin_out, cos_out);
                errors++;
            end else begin
                // Optional: Print latency for first few tests
                if (tests < 5) $display("Test %0d Passed. Latency: %0d cycles", tests, latency);
            end
            
            tests++;
            @(posedge clock); 
        end

        $display("Simulation Complete."); 
        $display("Tests: %0d, Errors: %0d", tests, errors);
        if (tests > 0) $display("Average Latency: %0.2f cycles", total_latency / tests);

        if (errors == 0) $display("SUCCESS: All tests passed.");
        else $display("FAILURE: %0d mismatches found.", errors);

        $fclose(rad_file);
        $fclose(sin_file);
        $fclose(cos_file);
        $finish;
    end

endmodule
