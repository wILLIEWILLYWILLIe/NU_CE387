
package cordic_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "cordic_global.sv"
    `include "cordic_transaction.sv"
    `include "cordic_sequence.sv"
    `include "cordic_monitor.sv"
    `include "cordic_driver.sv"
    `include "cordic_agent.sv"
    `include "cordic_scoreboard.sv"
    `include "cordic_env.sv"
    `include "cordic_test.sv"

endpackage
